module synth
(
    //io
)

    // body

endmodule