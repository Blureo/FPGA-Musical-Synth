module nco

// Waveform ROM
logic [15:0] waveform_rom [0:31];

// Waveform Slope ROM
logic [15:0] waveform_slope_rom [0:31];

endmodule